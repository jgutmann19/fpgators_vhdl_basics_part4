library ieee;
use ieee.std_logic_1164.all;

entity flip_flop is

end entity;